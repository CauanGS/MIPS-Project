library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ULA is
    Port (
        A, B : in std_logic_vector(31 downto 0);
        F : in std_logic_vector(2 downto 0);
        Y : out std_logic_vector(31 downto 0)
    );
end ULA;

architecture gate_level of ULA is
    signal BB : std_logic_vector(31 downto 0);
    signal S : std_logic_vector(31 downto 0);
begin

    process(A, B, F)
    begin
        if F(2) = '1' then
            BB <= B;
        else
            BB <= not B;
        end if;

        case F(1 downto 0) is
            when "00" =>
                Y <= A and B;
            when "01" =>
                Y <= A or B;
            when "11" =>
                S <= std_logic_vector(unsigned(A) + unsigned(not B) + 1);
                if F(0) = '1' then
                    if S(31) = '1' then
                        Y <= x"00000001";
                    else
                        Y <= x"00000000";
                    end if;
                else
                    Y <= S;
                end if;
            when others =>
                Y <= (others => '0');
        end case;
    end process;

end gate_level;
