library verilog;
use verilog.vl_types.all;
entity INST_MEM_vlg_vec_tst is
end INST_MEM_vlg_vec_tst;
